��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��㙂��c���љAtC�~�<ۼ���U�"�D��([z>��(gR�#���Zf�J�[���OE�X�#����z�3��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�`q�$&�[��!�2��T\!sw�����*o��]��0�P��%HJ�"�˽�Cd�}�Τ02��Yе
�#���R��_�3d#p�.5}�D����w4�>*A��%���:��dZ�x�cr��VQ6k�o�&�!=�@U�7��j�?�eG���8
��i.�-'� d���Y�|�O���ia9j!��wZ���4�d �Y�@<"������o���J}ƛY
��^�y��)߿�<�Փ?��؋�Mo�~��^r2"�:j!B��j>�p9�X��m��n����y����y>Q8�3sT��"����+�ɮ�@!�b�#U��ǫ�Rp�:n���հ���nz��,Ξ�Ӯ6�Ĕ,���w�{��=��f���Q�j�"檫5�j��b���L~#$���^�r�-����P�	�f�����g���l���*�J�w%)M�' �����!/ʦ�Qk4�;� �X�(�l{��+���_�
�lS��!�َ�(&��U�B{��4��.�n�ۼL��M/G�B��YГTK���M��7����%�,#��G/�8��s=�m�<�,\l�"M�u���6�۾YЖ�ܔ�{C���@�U����T�p������d��T���ԝ���w��@8D�s���4i�O�`.z/��q�C͠�'���ƣo=���a��X�Y����.���U`
n@i��-����#J��4��t5G)��D��'��h����c8C�f/Yls�X���9���>�?�R���P!��~�Y�[�=�@��%�����m�!s�d�E�s�{ |ö1�,\jmֽP.]�U����D&���P'K����I�2�e���c��B�]o �,-E��V��l�c����3{H�!D!r�w1�aE�wmڧ��?F��u��vrլ0�-��t�"��f�x�'D㩏�f'&��Ly�	��H�Lp��2����%	ׇ&��#&ti��EFeR	�����y;���Uv&w������� Ԁx�:��1�n.��Rg}��Q��;1@�D������އ�H�|jP*܃֟�AyΥ���}��r�@R�
�8��kh8��#%�k%�g��_�'�z)�վ@�,�>`T����h��zB�C���0�e*[o��Ao'cxZ�#���4i1�ӆ�����$�?�eZ�Z�F�B�?�k�e=�\�������3�x�6��,����%t��$g&��t�|�r�M�'�����C�e��3M���V�"�n�S7w+#�c�� ���������'�bƳ��B"�(E���?BM2��,�u÷ᴥ�U��U�?qw����ˤi.�@����i���� |��Hm��#]�7 �����;k�u�_����&Ĕ�B��[
��T�g�_~�b#:�TM*�3�]�e���՞$֊�u�:fn�2yn��+�̛�Śi��8E��p'|ө�i:a�v��TV�tu�B�¢����(��Άt(�,�}�t��1T���r�{��i��*�{����/ͤi��X�lBy�z_�up;1��b*��������L��N�`�xӤ{��s!�f�z��=�0MB}/�<�-YB�J����0ew�rx�����t�4�,��؟>�J���@[��$��nM{���F�����!fA��?#�V��������{u�x-z_6(Li ����d�K��Fz�I6\�&���v�}>��I�o�Ik�nz�d��ȃJ��S9� 2�z_�9Ҁ���d��"GM8	Ǟt�Ń�^�_ƽ)�o�~�Uv=װ s�<9$��c�'�թA����䟺6� �G1����15 9�
V�%p��^SZ�s�:[���>(Y���A��K����,�n��ch��h�!�m��+i���g��;c�E�z"\�������	[Vt�勗m��0(�� ��v>�h�̉O�R���QB�Ub�|��}���G����@�G��G�<W��X��^��3�>G�y�Zt�oc�S��R�*���&�S9S��%%v|������h:� ��Kj%��R��,9p��j���H����<<S�/?%�ƭis�P�I�S��s� �>��al���G���/�>�Hd{�,���rQ<��p�xJ�R�	Nw��'�\�Kp�����G�R׷����H��^h1�|<�M�&��AK�������IC=9��i��Y��xIԔҁ"���.�<K��F�_e�$d��ktΣ�`�/ϔ���oW?Y�CQN�k�wZk��Ȇs�if�fp�/�@���W�ܡz��5ĠC���;^}pN�껧������r������&��z��Ņ@/�ޑ(fO��Ć �	J.ANkw������t�G3ɻ��ߞ�xO<G��>����5ָ��V�����؏1`�?���[�'ra���Z-9Z���q���KaI�P�!bܔ�[OH!�D��2Q���M�����:���8��(ɟ0�����r��PK��TÄ��0{�tpJٸ.,ZYC�R��j�|�O!l�2F���[�K���x��!��TBfh%�
j�8I늎HHRO<糊 �Gɮ }ޣ��=�}��H��>�� ������~�$yJp2�ؼ��J��d�c���G�bL?6:�]k�2/�����,�Ǽ�B�(�ruI[h��8���dڇk���L+K��e�h��ݼ��_Q7��6��H
|�v}�Q�G� �ͦrh�E�cb���9�`skJ���f�܂Q1Ӡ���C����F�����w~�3�i�wA��i�x⾃4�'��^�{�s���ºY$���K�� �Bj��!��K�����x�}
�#n���=�V�=zv?6����!&*
��|�a��h!BK��M�����׹����K*΅\n���q��ֹq�T�xo��.�� p��1�zUwY6�|��?��쐻�Y���#uR?�l���v�����Y�!.�w��=f��L�y�t*���A�lM��_v�:wuh�&���e9JtNl�3�n)1
u�`a9��즐HhL�lYv���r���2I����F�푟���~v��d�������?�ϝ���P|�.�տ�ܟ�16��_vYڂ�La 	G��#�"�O���nమ�R���t��c"h���S��,d�]�-.]i���!.}��~{�hЊU�j�(�F/	�jU��_ś�)�h�$�>�/�l�ijݨ�S�xL�������bG��Y:VoB��}e�Z������D1��ݬ�Ɇ]�V��%�G�S����_Ԑ��b�S���������
���F��7,�l�l��;�S ���-b/,�[�T� �τfQjۙ,�ApIs��Mۡ��7���.��2T�3}%�YM@c�wb+��ƨ�R�x�ÏP�������\{)��35ƿj8�Dj��4� i���چ��ڞvgS��֯Li~������.��yYg(,.�2���F]��� ��}������cVq7��X��q��H��=��U.������44Qն#�`�v����:OX����j�)���n:|f��:�VR�zߢ��R�B�Q�j���WQK�*_'e6i?C���~�_�A�D�Ѱd�T�w�M�J����E�ע�l%3E��w�U����*m#x��!Z�{���|���ǮXP�����2���z�uf��/������F���/�a�q}*/���Dw��q� �|����N<$b��l�j7�YV�3'�:6xe�3G�pu�(�U#5A������ �&�������i�8�
�-�>���k�||�+(��g�<eb&�r�QVI3�Jĩ��s�-ᙀ��Q -�륗��>�ّᾐv��zr�~���@��C��M��R�2�v�ƾ䓎�C�^��g�Z�%b@��}�<,�d���YgŦ�ŁP��jO�S���D�z�nc�lӒ����}� _��]� Kp�|�����K�l^(A�
=5���J�)Q&��SZ��>�7���F�0����!^���b��7B'�F�.�h&d�r~�gG��:����W���t	�������w����|���N�HFs*\�6��e)���RP%GVl)v;�Pr����
�#�3Y��E���B��߹�rOKM�q�}e���:s����GeH|puÂ�CDJ?�%�G/�Xi�8�^���O���W��/�=�N;�v7��b���h���ػkô�M���)C�+�Z�T���ߴ�Re��A�*��<�S�^.٦����b�Ǝ�o��+�
�"A]o�$�ͅ�����2�9&�6�R��ә������a	����GNrc4�hp)4/�� l�y����E��E������a��״
c����쫥.]��GQ��ò�y�A��,�qn��[�