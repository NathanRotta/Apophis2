��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&r�F���ohC�*��}�o�r��t��W-T3.ϝ ]��K���k�U�����&�e\*$#��\�A����η�ɇk��%�ru�
��/@O�)���&���1�T m���������R���wfTS{����U�[J�� z�`������Α�%W�f[���U"*�BQ�`��8�O����꬛8,��9ҋr W%��+vF+���4|M8��k1�=꽧S�K�s4�ޣ�F�0��X�L���ֻ*LFh�ۼ��'|>'��	��hD���F��ݯu��'��_,[�����,�xEK��޽�#��G
QD"�l(e�A.�������8�P#5չ�̷�
�����)��7�m�Z�He�p�3��j{6W��o-��;���YШ�m�s]�{�Q4�̝I�b]X�̡߶��N\�d�\��E��'���P��c{��mo�՚n�G�d���5�)�D�4?�
F[�ʂ0�n|o*�DF%�E��LR��,�1d���).�u˪��%�SR��`���Q聨�hSR"��s�>!�����aS�p)I��b�i�mB
`��z�h����$��*�um�{��,� $�ePNR��v���}�Tn��w�G,V��M]����7�ߤ���1#�7[�j~��V�e�A�}�Aǅv&T�X"�6	YL.J�]FV�j��bo�q�r����z�g%=X��X����h�����,��Uf����}�{�=Z�j��Qa�����W�EMk�4�O}����7u`v��d[i�Y=X�� ��xnūH]P����������y�3��0�>Xi��i����Y}~��m^=��&i�G�o�f�K���S�|��+���Pe��i��fC�س- ��@S�! �`/�K�5�aك� �!�d2��i���A�G����7�R�7�Pʢ�5��図HQ)���	���ܘ0l���.�����Ɛ0��[2�j|��c=\�EX��������s7�~��s+�ڊ�Ȉ����C#e#Y}�O�n���e�z�O
IAo����T{�[8� r�O����f_����,m�6�G���`wj���;�h�^������@��A@��!Ɋ%���|6�A`�$I�ןN��>hh��:���}�ă��d\�����*�ӬÔ@��D�tݻq��[C�����V̤�T7!v�'I߃���մ
*���GI��Io&��$xefb�#o��gj�ߴCd�������BL��m��s𞖝9���2G#har-x�����x�jT�Vx��j�v�H����E��h��U\A<-�j-��n8b�I�e˕���8��u(����A��d��*M���"z[�(�~�ULT2��s$��aG���%��&�D�*o�:�d�v����uz��t�2	'Ty�=��F������%3����m=e^-��C~������ڥ����b6��*��ϗ����F���L�	�����ʤ�E�|Q��	+R��7��c��^��"��]���TZT��l��Zw��&���ʸ��ں�$�cd ��������nm0L���Q&�G�r)ۓ~���c�i�B&��u2�5h[D��X�����.}X��ތ���E����[,b�_|�z.	v��9�ۯ^�hY����c��s�7n�l\�-���@8��kB�`)���\2��Ξ��CE�z�V늑-Xf�Q	������k��w+L�E޻v|�R7�d��u�.��5�B���i��7|Dn�N \.r���FE�C�WK��ӗ��~��o�yk3X2��au�m�8a�NqF!�loÆD��$HY
�����<6��g[�s:�J?�	k���]a�N�Fwɻ���~+��u��Z�;���hYe�Cta���pEx�ɆR4�@��7?U-�
Re�����T�T(�k�I�܉��}�[�5IW�L�-���Do�dD1���U�Eym�Dq�d�?����FI�]Ŕ�Q�V?o��f$A��è���R�d��Q�^�#��)'�h2u�k���=��F�1��R���TZĠ2�,4Jͯ�qX�`�A���c��&�uDPBs���3H�/s���W~kH�a�Iz��Ij�MQu��:|P�C�\idĵ��5a>��:�?X<r3�ڙ6�=�v��Q@��g����nCOS�]O�(.0��}
���}+V������Q�"W�:��V�vJ��ަ�A޾��#�V���YƓ�@)m1@�ݜ���n2���5Vg)Y��z�IWg� a�
��3x=�m,�g�Oo�Ń'�*Kj�&��l�~�[p�u����f����Y�w0�z�Ph�>X"����$�1�.	RR�sXe��:���~�kA�������'xi2X��y�D%*�g×�E�?�ƻ(�h�VuZ���?�O�r,��|Su��@�[�C;8��Dw�"�}�QW��J�;{�'c3H�+H�^6�Q�LG�#���_����΂`��2KɚT&D�z�bzxѭ�P��F����H�z�hU�%�鋯�gl���IANK��n��!@OM�ֲ�$�t�O�wY6dU��q����xr/�Zk!UF�/3���d{��U��]�yr�+k���ĊT��ī8�qݐ�IFm���v�����Z]��uoM>�m;��p�j]7�Q$�}r�u.+���1*h6��T&�?e��"@Dbٟ-jN�y ������H�m.psL����g���c�M+4n�(q��T֬������B���!�� ��n���S��`&�:��L��t(��/SQ���9�j7�����HA�>�us9_z(����%��n�4Z
�Z�L,zQ%���b	{�!o s1sp\��Ϫ�2�{��FfU�ԠGT�;�J�8��|[׵���|�`)�|;���"j+p셚A������\~�Cx9� �2ё[�����t�'S�Qk(��v7n?i�k� �������:ڡ~��`?�)1!){�A���0���n�㻩W�8�,���_O�^�-a@�,��ٍA�"RU�G��>�l�Y8��	l�*��`���f
'��<�k=8Xe^4;ؘ�q"�9�,�1O����l	Z�B��JWpc����.��H��YД$�?�+9�iݗ��ڵC�_uٱ1�3�8
08��ه{TM[��)�`��<ga^��WBT��&͏Q��k�N�⤦.N\u�aH�G�Y�S]�����[���ĩ@{���$OiFÖpU�nJG���T(�Ϳ�/-�th\�ިA���tf�_��qW�8�������(�f>�������1v�\�G�����������7o!Ꚍ5���<�Du�K���r���j�\p^����J
��D��5Fnn�33:l�l��N�u�-��H�9�L[0��R�3@�f�5�KϨ�j�3���b<����9��v\=�3�C�d��?��[t�I�6b�f��L8_H��1��d�	 �섳q[o3[�G(hc򛈠�	�x�uBщ�ã)��vM6�@?̑��X|��u�.�9�#7�_��E$�|�sA�E�8U��ɦP&U>�R3J��%�=P}c�\?��M����T�=�`$H$���)`w�^�-4d��hHe�m��F�}��לů�RC=cwN�/��q:��֝���Җk7�w]��Xy��!*2�yC��GAjqX�ߦ~���&�Ԥ�^u��+l�3��n�T#�&�ؘ�6UG0q7�5���u��\�
q��`w�Qv�4)-~�ˀ�A0�kO��*��n������0��3�U,��@��X�2/� �BE�0��t���i�i�u%;�0όN�io�-�,�S��*&�+
��D�_�쉏^�Xp����8'$1F�הg}���:9�n��t^����t���
�G�z@]B�Sd�Z'$��C�	o��b]�Nn�@��'��)���S��6]C[_0�b��em�}X�鈾6�$']�����`��q�٘\ٵ���X�VNx�{���=��:`č���v�o�s��?$��uJ��E!yt�w��������d��cT��x�eb�������_�����Hr�j@B���*"�2 L�KX�&zc�ϫ�D���������Ȑ��{OC�b�!2�,f�U>R��H)�mVt6	��H]2
�@ȇ���6�d�'�:hRI
v��]N���e�Ӹp�}6�!;(N�dg����$�C� �R��ا"����$����~��q��X8@3\����ޠm��r�g�r�
6�X[>i#��\���پ.�p)_�k!�.��VM�Ƥ>F��*��;H͗��b���k=�̕ɱm*��u�U���}����S0�^R��J�I!~��
 ��="2��,0��3��*%����n��R��1:J uM��A����~�ϼ
X"Ǯ+ǔ�t�섭6�'�3���S#h����r��1�4MKy�����<�_b��p��i��h>�)�L��k�e%)�ë�vd�T����Ց�3$/�Hd�v�������i�nY~��EH��v�]���˧
�P�y%�'jYQ-A�:8s����������V������Tv�5;`�ΠR-p���N�ժ\W���\���H�	~Z+���g�tچX�#U	�[~#�+m�%ק����潢/�_��a8��|�f�gq~0>*ү��eQv��y�\>�E�� ���m��B�Y�Hp�zV��OV0�I�sߖ �o:��w�U�{��m��v�(����5r�Q���7]�8����?����W�w�dr�	K����Ȑ����P�^:�%�m��U�g��:��zhϏ%�ļ�ޗ��.�"��@�<��<��Q����}����K���r?��9y�HE}W֜�$b{��X	 ����j�_�~�s)k��^���6������m<�;̑�h�=>���OD���C�|j� φ��ĳծ���i^o��<_�n��׀DɎ���� ���I�C��� ���F����v:kw?��D�#3��G���%�/�ص^1������^�ڪU���O\+�]�5XMd˧D��[{Kkr�����~M?����7.��[1�^H����W`N���I�wc��*�Fk
���pM�}`K��A卣�+�Qs�F3�S
`AMY���e�
`b�_�����^2"�����H����<�Zh(=�3s�a2!Id�����7��)�ʄ]��mA��I��}��dfjXø!,.�˓��1���>�����	��p	7i�6�?h׆ΫcFEq?�Iy�@*����:�gۀ���1��
����t˜7�H��FI +���L�);�N7���H��2�:��v�6U6=I���[��˩�1֠���%[@ҿ�:�a(�D?��i�%� �f~�詁��_�C��m�c�Q\����m⫉�u$u�y"L�ʫ���F�⠴Ѩi�����![gּ�+3���x�<�.hC�=/^��O(�Xs.��c��B �~ T^?�Q���f�\���ƌ
�a7S6��©��O�3�]��Z��*�`��xo`b�.t��vA����	^�d�-��u��ɯ� 3���"O�������_IM7�D1��ʱ����ͳ��/�j�E\�5�� �ߥȳ����z����͛C�4���7�C{�t���p�����k���f�g(�Eo������;̡R����iN��<�$w�c���Ȥn�f�`	�oH7: �v-�����@=8�\(�k�,D�_�=�j^�=�&�;2�v�]d���ͻJ�=��@ôָ�z��T
��W�8��|+Y?���4�(}S�*,F2"(�y±�0�/�6G5�!� > m7���xȸn�7C��Do5�/JY�K�G"o^scl��G�z�B�!,���5�긢���4�W�3Z��\�4�2j�Q���B��Q*�;���wn�3�)ݧ@���w�:�n�n86�R���
Ѿ���c�F�^v8�ry�ėD�{�oN�"�8�4Њ�퇃��G�L86��h�~t���b��!��P!�*���I����v��eX5t3��/?^d�d�ٽ��8�j�N���e��Q�y[���8P���K� �4�	����\rju5�
4�S
��� ��$�v�7ʗ��U`d۾
�XY�,m��r�A��p/' �-�nJͅ�TT��rc����I1j�/i��/@Zb�Z
����X==�9�˕-{/&�ûE^�ؽ�feށE ������HNG_	�{�VEU�eA��#i�ո'3`��x�#�P��^M�{V$8
�e��+�a�����!eu:U��d1n��=uewe���\�Q'~Ne�����-�b�Np�1k�bZ�����,V��ǣ�5G��Ȭ3�V��H� ���s�	S�U����c��āN��]R��kP� ��e��;�:�8���<)n]'dڵ��m���7�Z�P�ʑ�;5��g����U���9��=����"D�oBܕ/������D��ж���A�`^q��3z�M�w�����$���D+�����$,�P[(ar����#�;7�v�Dc��:\��98�+�O+�cl���10ˊ�Pi���0���|�����uѻܒ@���)4�N��>����Wɕ����R}8�fȵQ5�G�1�,I��G�_��,u�&-�����_�!\7��o�vӇ\�1�b�P�'hn�&Z��x��"|�%i����T���% �N��բ���� 6�bЄp���_�s�*(oFv}q�<� #yA0� �3X�S����4b�9-���@8ş�c�%Ѿ���f^�&~�▾�]��ؓ?\��v��A�]]����X��M:��s#�E��)���gҷִ�!���<0`m��#����_t�!��L��L�/3t��}����__��p���
�a��grL�u���P{�C��kֱ~	�ݠ��^L�Tp>�3TTc�g
A��8D�y�{Q*.w��E9��j+�=�����ygU��D���/v[�ȩN퀋���#w��I@�'����2����w�ݽ�B��پԬ^Q��x�9�&Z��O�({������_U�4=�#C1�ʲf�4�2gWیc�P%��G	��ܛ�Tm�������{�{��7F�_�o��m�@0��`�SAG�J���P�%�{?D�8p:¡���qXT6?��8nυ���(!�7ͦ� eG��~ŋ�U�� +��0SDzp���^���o��&���j?�<v����?��u�2c�B�pCOH��%r̆D����=�+e?<�y��ΐknM6	uΎ��8�o�*�b�c�E:��J�Չ�Zў�,�� �5��@���AM��l��*_�O��ǳWߠx-cEj�N�BF)A~mYn�OĜ���n���)�d�nh���6���G���⬠���rĽ� y��u��M{���X�I��/�Q�`0��È�?�D�u?��e�Bi�?�ԭ���ɩ6��3r,��o[{��1�5��n`�ܿ(��r�V��8pӆ��Q�u>5�3-d1!⑒��Ҿ��h�����[�����n��P*%J;:���]���N��7��i����s�[����[v��z�����s@��O�B��d7~��M�2db�W8I/�_,�+!�m�x�����a�ի�X��7�4\�C�����Z����p�|��ԗS���
�g�Wc9L��R9�ɓ���	�i��!{fb7�(Ē,Ә-�R�a��1YA�7&�b:�G�o}R;9N�ǀ��5�_������k"rZA.0����W���JPh����E�$|��x6���-�Z�.s�� fCɟ�\��\� �8�w�n'��O�7_jv$�]d����f�?$��*��80v�2��&	w��
��ߣ��(�e�T��Q��:�9�􂊊O�U� N��e/�@i�49i��#騛���E_�D#��aӕ���M:!�672�����`�!+�\>P��\�y�nbh[���Ŷ�>ny,�vkH<j[�q��/��&ipX\ ��+��H��^�,�9����=�j脢L�{��,v����0�U�3z��� ���Ѯ���M̽����ZN�;�Hm==�\o�� <������xOL�Ӭ#Bj6/`�8���4���Ev��&y��c�ĩ3(L��I��hb��Vv�p��$��/����	nyF�������bNF^<5���Q?m