
`ifndef _macros_vh_
`define _macros_vh_
`define POW10(x) \
   (x == 0) ?  64'd1 : \
   (x == 1) ?  64'd10 : \
   (x == 2) ?  64'd100 : \
   (x == 3) ?  64'd1000 : \
   (x == 4) ?  64'd10000 : \
   (x == 5) ?  64'd100000 : \
   (x == 6) ?  64'd1000000 : \
   (x == 7) ?  64'd10000000 : \
   (x == 8) ?  64'd100000000 : \
   (x == 9) ?  64'd1000000000 : \
   (x == 10) ? 64'd10000000000 : \
   (x == 11) ? 64'd100000000000 : \
   (x == 12) ? 64'd1000000000000 : \
   (x == 13) ? 64'd10000000000000 : \
   (x == 14) ? 64'd100000000000000 : \
   (x == 15) ? 64'd1000000000000000 : \
   (x == 16) ? 64'd10000000000000000 : \
   (x == 17) ? 64'd100000000000000000 : \
   (x == 18) ? 64'd1000000000000000000 : \
   (x == 19) ? 64'd10000000000000000000 : \
   (x == 20) ? 64'd100000000000000000000 : \
   (x == 21) ? 64'd1000000000000000000000 : \
   (x == 22) ? 64'd10000000000000000000000 : \
   (x == 23) ? 64'd100000000000000000000000 : \
   (x == 24) ? 64'd1000000000000000000000000 : -1

`endif